module f3(a,b,c);
input [3:0]a,b,c;
wire [3:0]Y=a&b&c;
endmodule
